CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
68 C:\Users\phgi\~\Desktop\Arquivos\Programas\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 78 195 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
42711.2 0
0
13 Logic Switch~
5 77 157 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
42711.2 0
0
13 Logic Switch~
5 76 121 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
42711.2 0
0
7 Ground~
168 585 170 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3421 0 0
2
42711.2 0
0
4 LED~
171 498 106 0 2 2
10 6 2
0
0 0 864 90
4 LED0
-12 -21 16 -13
2 D4
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
8157 0 0
2
42711.2 0
0
4 LED~
171 438 105 0 2 2
10 7 2
0
0 0 864 90
4 LED0
-12 -21 16 -13
2 D3
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
5572 0 0
2
42711.2 0
0
4 LED~
171 379 103 0 2 2
10 8 2
0
0 0 864 90
4 LED0
-12 -21 16 -13
2 D2
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
8901 0 0
2
42711.2 0
0
4 LED~
171 326 104 0 2 2
10 9 2
0
0 0 864 90
4 LED0
-12 -21 16 -13
2 D1
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
7361 0 0
2
42711.2 0
0
4 4015
219 211 169 0 7 32
0 5 4 3 9 8 7 6
0
0 0 4848 0
4 4015
-14 -60 14 -52
3 U1A
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
65 %D [%16bi %8bi %1i %2i %3i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 9 6 5 4 3 10 7 9
6 5 4 3 10 15 1 14 13 12
11 2 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
4747 0 0
2
42711.2 0
0
11
1 3 3 0 0 4224 0 1 9 0 0 4
90 195
171 195
171 160
179 160
2 1 4 0 0 4224 0 9 2 0 0 4
179 142
98 142
98 157
89 157
1 1 5 0 0 4224 0 3 9 0 0 4
88 121
171 121
171 133
179 133
2 0 2 0 0 12416 0 8 0 0 7 4
339 105
367 105
367 136
585 136
2 0 2 0 0 0 0 7 0 0 7 4
392 104
426 104
426 128
585 128
2 0 2 0 0 0 0 6 0 0 7 2
451 106
585 107
2 1 2 0 0 0 0 5 4 0 0 3
511 107
585 107
585 164
7 1 6 0 0 4224 0 9 5 0 0 4
243 133
482 133
482 107
491 107
6 1 7 0 0 4224 0 9 6 0 0 4
243 142
422 142
422 106
431 106
5 1 8 0 0 4224 0 9 7 0 0 4
243 151
363 151
363 104
372 104
4 1 9 0 0 4224 0 9 8 0 0 4
243 160
310 160
310 105
319 105
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
